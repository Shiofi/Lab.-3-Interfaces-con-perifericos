`timescale 1ns / 1ps

module tb_UART_top(

);
endmodule