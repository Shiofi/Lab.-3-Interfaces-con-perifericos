`timescale 1ns / 1ps

module ControlReg (
    input logic clk, rst,
    input logic [31:0] IN1,
    input logic [31:0] IN2,
    input logic WR1,
    input logic WR2,
    output logic out
);


endmodule